signal sigA, sigB, sigC, sigN : 6;



sigA <= do something else;
p <= do something;