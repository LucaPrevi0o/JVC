signal sigA, sigB, sigC, sigN: std_logic_vector(2 to 4);
signal a, sgbgbeh, c, d, e, f: bit;
